`ifndef clocks_vh
`define clocks_vh

`define CLK_1X_WIDESCREEN 16875000
`define CLK_1X_STANDARD 12587500
`define CLK_2X_WIDESCREEN 33750000
`define CLK_2X_STANDARD 25175000


`endif

